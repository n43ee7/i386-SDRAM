module PLLVCO2 (
	input CLK,
	output READY,
	output CLKOUT

);

endmodule 